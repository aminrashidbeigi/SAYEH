library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity tan_co is
	port (
	input : in std_logic_vector(15 DOWNTO 0);
	output : out std_logic_vector(15 DOWNTO 0)
	);
end entity ;

architecture rtl of tan_co is

begin
	output <=
			"0000000000000000" when input = "0000000000000000" else
			"0000000000000000" when input = "0000000000000001" else
			"0000000000000000" when input = "0000000000000010" else
			"0000000000000000" when input = "0000000000000011" else
			"0000000000000000" when input = "0000000000000100" else
			"0000000000000000" when input = "0000000000000101" else
			"0000000000000001" when input = "0000000000000110" else
			"0000000000000001" when input = "0000000000000111" else
			"0000000000000001" when input = "0000000000001000" else
			"0000000000000001" when input = "0000000000001001" else
			"0000000000000001" when input = "0000000000001010" else
			"0000000000000001" when input = "0000000000001011" else
			"0000000000000010" when input = "0000000000001100" else
			"0000000000000010" when input = "0000000000001101" else
			"0000000000000010" when input = "0000000000001110" else
			"0000000000000010" when input = "0000000000001111" else
			"0000000000000010" when input = "0000000000010000" else
			"0000000000000011" when input = "0000000000010001" else
			"0000000000000011" when input = "0000000000010010" else
			"0000000000000011" when input = "0000000000010011" else
			"0000000000000011" when input = "0000000000010100" else
			"0000000000000011" when input = "0000000000010101" else
			"0000000000000100" when input = "0000000000010110" else
			"0000000000000100" when input = "0000000000010111" else
			"0000000000000100" when input = "0000000000011000" else
			"0000000000000100" when input = "0000000000011001" else
			"0000000000000100" when input = "0000000000011010" else
			"0000000000000101" when input = "0000000000011011" else
			"0000000000000101" when input = "0000000000011100" else
			"0000000000000101" when input = "0000000000011101" else
			"0000000000000101" when input = "0000000000011110" else
			"0000000000000110" when input = "0000000000011111" else
			"0000000000000110" when input = "0000000000100000" else
			"0000000000000110" when input = "0000000000100001" else
			"0000000000000110" when input = "0000000000100010" else
			"0000000000000111" when input = "0000000000100011" else
			"0000000000000111" when input = "0000000000100100" else
			"0000000000000111" when input = "0000000000100101" else
			"0000000000000111" when input = "0000000000100110" else
			"0000000000001000" when input = "0000000000100111" else
			"0000000000001000" when input = "0000000000101000" else
			"0000000000001000" when input = "0000000000101001" else
			"0000000000001001" when input = "0000000000101010" else
			"0000000000001001" when input = "0000000000101011" else
			"0000000000001001" when input = "0000000000101100" else
			"0000000000001001" when input = "0000000000101101" else
			"0000000000001010" when input = "0000000000101110" else
			"0000000000001010" when input = "0000000000101111" else
			"0000000000001011" when input = "0000000000110000" else
			"0000000000001011" when input = "0000000000110001" else
			"0000000000001011" when input = "0000000000110010" else
			"0000000000001100" when input = "0000000000110011" else
			"0000000000001100" when input = "0000000000110100" else
			"0000000000001101" when input = "0000000000110101" else
			"0000000000001101" when input = "0000000000110110" else
			"0000000000001110" when input = "0000000000110111" else
			"0000000000001110" when input = "0000000000111000" else
			"0000000000001111" when input = "0000000000111001" else
			"0000000000010000" when input = "0000000000111010" else
			"0000000000010000" when input = "0000000000111011" else
			"0000000000010001" when input = "0000000000111100" else
			"0000000000010010" when input = "0000000000111101" else
			"0000000000010010" when input = "0000000000111110" else
			"0000000000010011" when input = "0000000000111111" else
			"0000000000010100" when input = "0000000001000000" else
			"0000000000010101" when input = "0000000001000001" else
			"0000000000010110" when input = "0000000001000010" else
			"0000000000010111" when input = "0000000001000011" else
			"0000000000011000" when input = "0000000001000100" else
			"0000000000011010" when input = "0000000001000101" else
			"0000000000011011" when input = "0000000001000110" else
			"0000000000011101" when input = "0000000001000111" else
			"0000000000011110" when input = "0000000001001000" else
			"0000000000100000" when input = "0000000001001001" else
			"0000000000100010" when input = "0000000001001010" else
			"0000000000100101" when input = "0000000001001011" else
			"0000000000101000" when input = "0000000001001100" else
			"0000000000101011" when input = "0000000001001101" else
			"0000000000101111" when input = "0000000001001110" else
			"0000000000110011" when input = "0000000001001111" else
			"0000000000111000" when input = "0000000001010000" else
			"0000000000111111" when input = "0000000001010001" else
			"0000000001000111" when input = "0000000001010010" else
			"0000000001010001" when input = "0000000001010011" else
			"0000000001011111" when input = "0000000001010100" else
			"0000000001110010" when input = "0000000001010101" else
			"0000000010001110" when input = "0000000001010110" else
			"0000000010111110" when input = "0000000001010111" else
			"0000000100011101" when input = "0000000001011000" else
			"0000001000111011" when input = "0000000001011001" else
			"0100101100110001" when input = "0000000001011010" else
			"1111110111000010" when input = "0000000001011011" else
			"1111111011100010" when input = "0000000001011100" else
			"1111111101000010" when input = "0000000001011101" else
			"1111111101110001" when input = "0000000001011110" else
			"1111111110001110" when input = "0000000001011111" else
			"1111111110100001" when input = "0000000001100000" else
			"1111111110101111" when input = "0000000001100001" else
			"1111111110111001" when input = "0000000001100010" else
			"1111111111000001" when input = "0000000001100011" else
			"1111111111001000" when input = "0000000001100100" else
			"1111111111001101" when input = "0000000001100101" else
			"1111111111010001" when input = "0000000001100110" else
			"1111111111010101" when input = "0000000001100111" else
			"1111111111011000" when input = "0000000001101000" else
			"1111111111011011" when input = "0000000001101001" else
			"1111111111011110" when input = "0000000001101010" else
			"1111111111100000" when input = "0000000001101011" else
			"1111111111100010" when input = "0000000001101100" else
			"1111111111100011" when input = "0000000001101101" else
			"1111111111100101" when input = "0000000001101110" else
			"1111111111100110" when input = "0000000001101111" else
			"1111111111101000" when input = "0000000001110000" else
			"1111111111101001" when input = "0000000001110001" else
			"1111111111101010" when input = "0000000001110010" else
			"1111111111101011" when input = "0000000001110011" else
			"1111111111101100" when input = "0000000001110100" else
			"1111111111101101" when input = "0000000001110101" else
			"1111111111101110" when input = "0000000001110110" else
			"1111111111101110" when input = "0000000001110111" else
			"1111111111101111" when input = "0000000001111000" else
			"1111111111110000" when input = "0000000001111001" else
			"1111111111110000" when input = "0000000001111010" else
			"1111111111110001" when input = "0000000001111011" else
			"1111111111110010" when input = "0000000001111100" else
			"1111111111110010" when input = "0000000001111101" else
			"1111111111110011" when input = "0000000001111110" else
			"1111111111110011" when input = "0000000001111111" else
			"1111111111110100" when input = "0000000010000000" else
			"1111111111110100" when input = "0000000010000001" else
			"1111111111110101" when input = "0000000010000010" else
			"1111111111110101" when input = "0000000010000011" else
			"1111111111110101" when input = "0000000010000100" else
			"1111111111110110" when input = "0000000010000101" else
			"1111111111110110" when input = "0000000010000110" else
			"1111111111110110" when input = "0000000010000111" else
			"1111111111110111" when input = "0000000010001000" else
			"1111111111110111" when input = "0000000010001001" else
			"1111111111110111" when input = "0000000010001010" else
			"1111111111111000" when input = "0000000010001011" else
			"1111111111111000" when input = "0000000010001100" else
			"1111111111111000" when input = "0000000010001101" else
			"1111111111111001" when input = "0000000010001110" else
			"1111111111111001" when input = "0000000010001111" else
			"1111111111111001" when input = "0000000010010000" else
			"1111111111111001" when input = "0000000010010001" else
			"1111111111111010" when input = "0000000010010010" else
			"1111111111111010" when input = "0000000010010011" else
			"1111111111111010" when input = "0000000010010100" else
			"1111111111111010" when input = "0000000010010101" else
			"1111111111111011" when input = "0000000010010110" else
			"1111111111111011" when input = "0000000010010111" else
			"1111111111111011" when input = "0000000010011000" else
			"1111111111111011" when input = "0000000010011001" else
			"1111111111111100" when input = "0000000010011010" else
			"1111111111111100" when input = "0000000010011011" else
			"1111111111111100" when input = "0000000010011100" else
			"1111111111111100" when input = "0000000010011101" else
			"1111111111111100" when input = "0000000010011110" else
			"1111111111111101" when input = "0000000010011111" else
			"1111111111111101" when input = "0000000010100000" else
			"1111111111111101" when input = "0000000010100001" else
			"1111111111111101" when input = "0000000010100010" else
			"1111111111111101" when input = "0000000010100011" else
			"1111111111111110" when input = "0000000010100100" else
			"1111111111111110" when input = "0000000010100101" else
			"1111111111111110" when input = "0000000010100110" else
			"1111111111111110" when input = "0000000010100111" else
			"1111111111111110" when input = "0000000010101000" else
			"1111111111111111" when input = "0000000010101001" else
			"1111111111111111" when input = "0000000010101010" else
			"1111111111111111" when input = "0000000010101011" else
			"1111111111111111" when input = "0000000010101100" else
			"1111111111111111" when input = "0000000010101101" else
			"1111111111111111" when input = "0000000010101110" else
			"0000000000000000" when input = "0000000010101111" else
			"0000000000000000" when input = "0000000010110000" else
			"0000000000000000" when input = "0000000010110001" else
			"0000000000000000" when input = "0000000010110010" else
			"0000000000000000" when input = "0000000010110011" else
			"0000000000000000" when input = "0000000010110100" else
			"0000000000000000" when input = "0000000010110101" else
			"0000000000000000" when input = "0000000010110110" else
			"0000000000000000" when input = "0000000010110111" else
			"0000000000000000" when input = "0000000010111000" else
			"0000000000000000" when input = "0000000010111001" else
			"0000000000000001" when input = "0000000010111010" else
			"0000000000000001" when input = "0000000010111011" else
			"0000000000000001" when input = "0000000010111100" else
			"0000000000000001" when input = "0000000010111101" else
			"0000000000000001" when input = "0000000010111110" else
			"0000000000000001" when input = "0000000010111111" else
			"0000000000000010" when input = "0000000011000000" else
			"0000000000000010" when input = "0000000011000001" else
			"0000000000000010" when input = "0000000011000010" else
			"0000000000000010" when input = "0000000011000011" else
			"0000000000000010" when input = "0000000011000100" else
			"0000000000000011" when input = "0000000011000101" else
			"0000000000000011" when input = "0000000011000110" else
			"0000000000000011" when input = "0000000011000111" else
			"0000000000000011" when input = "0000000011001000" else
			"0000000000000011" when input = "0000000011001001" else
			"0000000000000100" when input = "0000000011001010" else
			"0000000000000100" when input = "0000000011001011" else
			"0000000000000100" when input = "0000000011001100" else
			"0000000000000100" when input = "0000000011001101" else
			"0000000000000100" when input = "0000000011001110" else
			"0000000000000101" when input = "0000000011001111" else
			"0000000000000101" when input = "0000000011010000" else
			"0000000000000101" when input = "0000000011010001" else
			"0000000000000101" when input = "0000000011010010" else
			"0000000000000110" when input = "0000000011010011" else
			"0000000000000110" when input = "0000000011010100" else
			"0000000000000110" when input = "0000000011010101" else
			"0000000000000110" when input = "0000000011010110" else
			"0000000000000111" when input = "0000000011010111" else
			"0000000000000111" when input = "0000000011011000" else
			"0000000000000111" when input = "0000000011011001" else
			"0000000000000111" when input = "0000000011011010" else
			"0000000000001000" when input = "0000000011011011" else
			"0000000000001000" when input = "0000000011011100" else
			"0000000000001000" when input = "0000000011011101" else
			"0000000000001001" when input = "0000000011011110" else
			"0000000000001001" when input = "0000000011011111" else
			"0000000000001001" when input = "0000000011100000" else
			"0000000000001001" when input = "0000000011100001" else
			"0000000000001010" when input = "0000000011100010" else
			"0000000000001010" when input = "0000000011100011" else
			"0000000000001011" when input = "0000000011100100" else
			"0000000000001011" when input = "0000000011100101" else
			"0000000000001011" when input = "0000000011100110" else
			"0000000000001100" when input = "0000000011100111" else
			"0000000000001100" when input = "0000000011101000" else
			"0000000000001101" when input = "0000000011101001" else
			"0000000000001101" when input = "0000000011101010" else
			"0000000000001110" when input = "0000000011101011" else
			"0000000000001110" when input = "0000000011101100" else
			"0000000000001111" when input = "0000000011101101" else
			"0000000000001111" when input = "0000000011101110" else
			"0000000000010000" when input = "0000000011101111" else
			"0000000000010001" when input = "0000000011110000" else
			"0000000000010010" when input = "0000000011110001" else
			"0000000000010010" when input = "0000000011110010" else
			"0000000000010011" when input = "0000000011110011" else
			"0000000000010100" when input = "0000000011110100" else
			"0000000000010101" when input = "0000000011110101" else
			"0000000000010110" when input = "0000000011110110" else
			"0000000000010111" when input = "0000000011110111" else
			"0000000000011000" when input = "0000000011111000" else
			"0000000000011010" when input = "0000000011111001" else
			"0000000000011011" when input = "0000000011111010" else
			"0000000000011101" when input = "0000000011111011" else
			"0000000000011110" when input = "0000000011111100" else
			"0000000000100000" when input = "0000000011111101" else
			"0000000000100010" when input = "0000000011111110" else
			"0000000000100101" when input = "0000000011111111" else
			"0000000000101000" when input = "0000000100000000" else
			"0000000000101011" when input = "0000000100000001" else
			"0000000000101111" when input = "0000000100000010" else
			"0000000000110011" when input = "0000000100000011" else
			"0000000000111000" when input = "0000000100000100" else
			"0000000000111111" when input = "0000000100000101" else
			"0000000001000111" when input = "0000000100000110" else
			"0000000001010001" when input = "0000000100000111" else
			"0000000001011111" when input = "0000000100001000" else
			"0000000001110010" when input = "0000000100001001" else
			"0000000010001110" when input = "0000000100001010" else
			"0000000010111110" when input = "0000000100001011" else
			"0000000100011101" when input = "0000000100001100" else
			"0000001000111000" when input = "0000000100001101" else
			"0001100100010000" when input = "0000000100001110" else
			"1111110110111111" when input = "0000000100001111" else
			"1111111011100001" when input = "0000000100010000" else
			"1111111101000001" when input = "0000000100010001" else
			"1111111101110001" when input = "0000000100010010" else
			"1111111110001110" when input = "0000000100010011" else
			"1111111110100001" when input = "0000000100010100" else
			"1111111110101111" when input = "0000000100010101" else
			"1111111110111001" when input = "0000000100010110" else
			"1111111111000001" when input = "0000000100010111" else
			"1111111111001000" when input = "0000000100011000" else
			"1111111111001101" when input = "0000000100011001" else
			"1111111111010001" when input = "0000000100011010" else
			"1111111111010101" when input = "0000000100011011" else
			"1111111111011000" when input = "0000000100011100" else
			"1111111111011011" when input = "0000000100011101" else
			"1111111111011110" when input = "0000000100011110" else
			"1111111111100000" when input = "0000000100011111" else
			"1111111111100010" when input = "0000000100100000" else
			"1111111111100011" when input = "0000000100100001" else
			"1111111111100101" when input = "0000000100100010" else
			"1111111111100110" when input = "0000000100100011" else
			"1111111111101000" when input = "0000000100100100" else
			"1111111111101001" when input = "0000000100100101" else
			"1111111111101010" when input = "0000000100100110" else
			"1111111111101011" when input = "0000000100100111" else
			"1111111111101100" when input = "0000000100101000" else
			"1111111111101101" when input = "0000000100101001" else
			"1111111111101110" when input = "0000000100101010" else
			"1111111111101110" when input = "0000000100101011" else
			"1111111111101111" when input = "0000000100101100" else
			"1111111111110000" when input = "0000000100101101" else
			"1111111111110000" when input = "0000000100101110" else
			"1111111111110001" when input = "0000000100101111" else
			"1111111111110010" when input = "0000000100110000" else
			"1111111111110010" when input = "0000000100110001" else
			"1111111111110011" when input = "0000000100110010" else
			"1111111111110011" when input = "0000000100110011" else
			"1111111111110100" when input = "0000000100110100" else
			"1111111111110100" when input = "0000000100110101" else
			"1111111111110101" when input = "0000000100110110" else
			"1111111111110101" when input = "0000000100110111" else
			"1111111111110101" when input = "0000000100111000" else
			"1111111111110110" when input = "0000000100111001" else
			"1111111111110110" when input = "0000000100111010" else
			"1111111111110110" when input = "0000000100111011" else
			"1111111111110111" when input = "0000000100111100" else
			"1111111111110111" when input = "0000000100111101" else
			"1111111111110111" when input = "0000000100111110" else
			"1111111111111000" when input = "0000000100111111" else
			"1111111111111000" when input = "0000000101000000" else
			"1111111111111000" when input = "0000000101000001" else
			"1111111111111001" when input = "0000000101000010" else
			"1111111111111001" when input = "0000000101000011" else
			"1111111111111001" when input = "0000000101000100" else
			"1111111111111001" when input = "0000000101000101" else
			"1111111111111010" when input = "0000000101000110" else
			"1111111111111010" when input = "0000000101000111" else
			"1111111111111010" when input = "0000000101001000" else
			"1111111111111010" when input = "0000000101001001" else
			"1111111111111011" when input = "0000000101001010" else
			"1111111111111011" when input = "0000000101001011" else
			"1111111111111011" when input = "0000000101001100" else
			"1111111111111011" when input = "0000000101001101" else
			"1111111111111100" when input = "0000000101001110" else
			"1111111111111100" when input = "0000000101001111" else
			"1111111111111100" when input = "0000000101010000" else
			"1111111111111100" when input = "0000000101010001" else
			"1111111111111100" when input = "0000000101010010" else
			"1111111111111101" when input = "0000000101010011" else
			"1111111111111101" when input = "0000000101010100" else
			"1111111111111101" when input = "0000000101010101" else
			"1111111111111101" when input = "0000000101010110" else
			"1111111111111101" when input = "0000000101010111" else
			"1111111111111110" when input = "0000000101011000" else
			"1111111111111110" when input = "0000000101011001" else
			"1111111111111110" when input = "0000000101011010" else
			"1111111111111110" when input = "0000000101011011" else
			"1111111111111110" when input = "0000000101011100" else
			"1111111111111111" when input = "0000000101011101" else
			"1111111111111111" when input = "0000000101011110" else
			"1111111111111111" when input = "0000000101011111" else
			"1111111111111111" when input = "0000000101100000" else
			"1111111111111111" when input = "0000000101100001" else
			"1111111111111111" when input = "0000000101100010" else
			"0000000000000000" when input = "0000000101100011" else
			"0000000000000000" when input = "0000000101100100" else
			"0000000000000000" when input = "0000000101100101" else
			"0000000000000000" when input = "0000000101100110" else
			"0000000000000000" when input = "0000000101100111" else
			"0000000000000000" when input = "0000000101101000" else
			"XXXXXXXXXXXXXXXX";
end architecture;
