library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity cos_co is
	port (
	input : in std_logic_vector(15 DOWNTO 0);
	output : out std_logic_vector(15 DOWNTO 0)
	);
end cos_co;

architecture rtl of cos_co is
begin
	output <=
			"0000001111101000" when input = "0000000000000000" else
			"0000001111100111" when input = "0000000000000001" else
			"0000001111100111" when input = "0000000000000010" else
			"0000001111100110" when input = "0000000000000011" else
			"0000001111100101" when input = "0000000000000100" else
			"0000001111100100" when input = "0000000000000101" else
			"0000001111100010" when input = "0000000000000110" else
			"0000001111100000" when input = "0000000000000111" else
			"0000001111011110" when input = "0000000000001000" else
			"0000001111011011" when input = "0000000000001001" else
			"0000001111011000" when input = "0000000000001010" else
			"0000001111010101" when input = "0000000000001011" else
			"0000001111010010" when input = "0000000000001100" else
			"0000001111001110" when input = "0000000000001101" else
			"0000001111001010" when input = "0000000000001110" else
			"0000001111000101" when input = "0000000000001111" else
			"0000001111000001" when input = "0000000000010000" else
			"0000001110111100" when input = "0000000000010001" else
			"0000001110110111" when input = "0000000000010010" else
			"0000001110110001" when input = "0000000000010011" else
			"0000001110101011" when input = "0000000000010100" else
			"0000001110100101" when input = "0000000000010101" else
			"0000001110011111" when input = "0000000000010110" else
			"0000001110011000" when input = "0000000000010111" else
			"0000001110010001" when input = "0000000000011000" else
			"0000001110001010" when input = "0000000000011001" else
			"0000001110000010" when input = "0000000000011010" else
			"0000001101111011" when input = "0000000000011011" else
			"0000001101110010" when input = "0000000000011100" else
			"0000001101101010" when input = "0000000000011101" else
			"0000001101100010" when input = "0000000000011110" else
			"0000001101011001" when input = "0000000000011111" else
			"0000001101010000" when input = "0000000000100000" else
			"0000001101000110" when input = "0000000000100001" else
			"0000001100111101" when input = "0000000000100010" else
			"0000001100110011" when input = "0000000000100011" else
			"0000001100101001" when input = "0000000000100100" else
			"0000001100011110" when input = "0000000000100101" else
			"0000001100010100" when input = "0000000000100110" else
			"0000001100001001" when input = "0000000000100111" else
			"0000001011111110" when input = "0000000000101000" else
			"0000001011110010" when input = "0000000000101001" else
			"0000001011100111" when input = "0000000000101010" else
			"0000001011011011" when input = "0000000000101011" else
			"0000001011001111" when input = "0000000000101100" else
			"0000001011000011" when input = "0000000000101101" else
			"0000001010110110" when input = "0000000000101110" else
			"0000001010101010" when input = "0000000000101111" else
			"0000001010011101" when input = "0000000000110000" else
			"0000001010010000" when input = "0000000000110001" else
			"0000001010000010" when input = "0000000000110010" else
			"0000001001110101" when input = "0000000000110011" else
			"0000001001100111" when input = "0000000000110100" else
			"0000001001011001" when input = "0000000000110101" else
			"0000001001001011" when input = "0000000000110110" else
			"0000001000111101" when input = "0000000000110111" else
			"0000001000101111" when input = "0000000000111000" else
			"0000001000100000" when input = "0000000000111001" else
			"0000001000010001" when input = "0000000000111010" else
			"0000001000000011" when input = "0000000000111011" else
			"0000000111110100" when input = "0000000000111100" else
			"0000000111100100" when input = "0000000000111101" else
			"0000000111010101" when input = "0000000000111110" else
			"0000000111000110" when input = "0000000000111111" else
			"0000000110110110" when input = "0000000001000000" else
			"0000000110100110" when input = "0000000001000001" else
			"0000000110010110" when input = "0000000001000010" else
			"0000000110000110" when input = "0000000001000011" else
			"0000000101110110" when input = "0000000001000100" else
			"0000000101100110" when input = "0000000001000101" else
			"0000000101010110" when input = "0000000001000110" else
			"0000000101000101" when input = "0000000001000111" else
			"0000000100110101" when input = "0000000001001000" else
			"0000000100100100" when input = "0000000001001001" else
			"0000000100010011" when input = "0000000001001010" else
			"0000000100000010" when input = "0000000001001011" else
			"0000000011110001" when input = "0000000001001100" else
			"0000000011100000" when input = "0000000001001101" else
			"0000000011001111" when input = "0000000001001110" else
			"0000000010111110" when input = "0000000001001111" else
			"0000000010101101" when input = "0000000001010000" else
			"0000000010011100" when input = "0000000001010001" else
			"0000000010001011" when input = "0000000001010010" else
			"0000000001111001" when input = "0000000001010011" else
			"0000000001101000" when input = "0000000001010100" else
			"0000000001010111" when input = "0000000001010101" else
			"0000000001000101" when input = "0000000001010110" else
			"0000000000110100" when input = "0000000001010111" else
			"0000000000100010" when input = "0000000001011000" else
			"0000000000010001" when input = "0000000001011001" else
			"0000000000000000" when input = "0000000001011010" else
			"1111111111101111" when input = "0000000001011011" else
			"1111111111011110" when input = "0000000001011100" else
			"1111111111001100" when input = "0000000001011101" else
			"1111111110111011" when input = "0000000001011110" else
			"1111111110101001" when input = "0000000001011111" else
			"1111111110011000" when input = "0000000001100000" else
			"1111111110000111" when input = "0000000001100001" else
			"1111111101110101" when input = "0000000001100010" else
			"1111111101100100" when input = "0000000001100011" else
			"1111111101010011" when input = "0000000001100100" else
			"1111111101000010" when input = "0000000001100101" else
			"1111111100110001" when input = "0000000001100110" else
			"1111111100100000" when input = "0000000001100111" else
			"1111111100001111" when input = "0000000001101000" else
			"1111111011111110" when input = "0000000001101001" else
			"1111111011101101" when input = "0000000001101010" else
			"1111111011011100" when input = "0000000001101011" else
			"1111111011001100" when input = "0000000001101100" else
			"1111111010111011" when input = "0000000001101101" else
			"1111111010101011" when input = "0000000001101110" else
			"1111111010011010" when input = "0000000001101111" else
			"1111111010001010" when input = "0000000001110000" else
			"1111111001111010" when input = "0000000001110001" else
			"1111111001101010" when input = "0000000001110010" else
			"1111111001011010" when input = "0000000001110011" else
			"1111111001001010" when input = "0000000001110100" else
			"1111111000111011" when input = "0000000001110101" else
			"1111111000101011" when input = "0000000001110110" else
			"1111111000011100" when input = "0000000001110111" else
			"1111111000001101" when input = "0000000001111000" else
			"1111110111111110" when input = "0000000001111001" else
			"1111110111101111" when input = "0000000001111010" else
			"1111110111100000" when input = "0000000001111011" else
			"1111110111010001" when input = "0000000001111100" else
			"1111110111000011" when input = "0000000001111101" else
			"1111110110110101" when input = "0000000001111110" else
			"1111110110100111" when input = "0000000001111111" else
			"1111110110011001" when input = "0000000010000000" else
			"1111110110001011" when input = "0000000010000001" else
			"1111110101111110" when input = "0000000010000010" else
			"1111110101110000" when input = "0000000010000011" else
			"1111110101100011" when input = "0000000010000100" else
			"1111110101010111" when input = "0000000010000101" else
			"1111110101001010" when input = "0000000010000110" else
			"1111110100111101" when input = "0000000010000111" else
			"1111110100110001" when input = "0000000010001000" else
			"1111110100100101" when input = "0000000010001001" else
			"1111110100011001" when input = "0000000010001010" else
			"1111110100001110" when input = "0000000010001011" else
			"1111110100000011" when input = "0000000010001100" else
			"1111110011110111" when input = "0000000010001101" else
			"1111110011101101" when input = "0000000010001110" else
			"1111110011100010" when input = "0000000010001111" else
			"1111110011011000" when input = "0000000010010000" else
			"1111110011001101" when input = "0000000010010001" else
			"1111110011000100" when input = "0000000010010010" else
			"1111110010111010" when input = "0000000010010011" else
			"1111110010110000" when input = "0000000010010100" else
			"1111110010100111" when input = "0000000010010101" else
			"1111110010011111" when input = "0000000010010110" else
			"1111110010010110" when input = "0000000010010111" else
			"1111110010001110" when input = "0000000010011000" else
			"1111110010000110" when input = "0000000010011001" else
			"1111110001111110" when input = "0000000010011010" else
			"1111110001110110" when input = "0000000010011011" else
			"1111110001101111" when input = "0000000010011100" else
			"1111110001101000" when input = "0000000010011101" else
			"1111110001100001" when input = "0000000010011110" else
			"1111110001011011" when input = "0000000010011111" else
			"1111110001010101" when input = "0000000010100000" else
			"1111110001001111" when input = "0000000010100001" else
			"1111110001001001" when input = "0000000010100010" else
			"1111110001000100" when input = "0000000010100011" else
			"1111110000111111" when input = "0000000010100100" else
			"1111110000111011" when input = "0000000010100101" else
			"1111110000110110" when input = "0000000010100110" else
			"1111110000110010" when input = "0000000010100111" else
			"1111110000101110" when input = "0000000010101000" else
			"1111110000101011" when input = "0000000010101001" else
			"1111110000101000" when input = "0000000010101010" else
			"1111110000100101" when input = "0000000010101011" else
			"1111110000100010" when input = "0000000010101100" else
			"1111110000100000" when input = "0000000010101101" else
			"1111110000011110" when input = "0000000010101110" else
			"1111110000011100" when input = "0000000010101111" else
			"1111110000011011" when input = "0000000010110000" else
			"1111110000011010" when input = "0000000010110001" else
			"1111110000011001" when input = "0000000010110010" else
			"1111110000011001" when input = "0000000010110011" else
			"1111110000011001" when input = "0000000010110100" else
			"1111110000011001" when input = "0000000010110101" else
			"1111110000011001" when input = "0000000010110110" else
			"1111110000011010" when input = "0000000010110111" else
			"1111110000011011" when input = "0000000010111000" else
			"1111110000011100" when input = "0000000010111001" else
			"1111110000011110" when input = "0000000010111010" else
			"1111110000100000" when input = "0000000010111011" else
			"1111110000100010" when input = "0000000010111100" else
			"1111110000100101" when input = "0000000010111101" else
			"1111110000101000" when input = "0000000010111110" else
			"1111110000101011" when input = "0000000010111111" else
			"1111110000101110" when input = "0000000011000000" else
			"1111110000110010" when input = "0000000011000001" else
			"1111110000110110" when input = "0000000011000010" else
			"1111110000111011" when input = "0000000011000011" else
			"1111110000111111" when input = "0000000011000100" else
			"1111110001000100" when input = "0000000011000101" else
			"1111110001001001" when input = "0000000011000110" else
			"1111110001001111" when input = "0000000011000111" else
			"1111110001010101" when input = "0000000011001000" else
			"1111110001011011" when input = "0000000011001001" else
			"1111110001100001" when input = "0000000011001010" else
			"1111110001101000" when input = "0000000011001011" else
			"1111110001101111" when input = "0000000011001100" else
			"1111110001110110" when input = "0000000011001101" else
			"1111110001111110" when input = "0000000011001110" else
			"1111110010000101" when input = "0000000011001111" else
			"1111110010001110" when input = "0000000011010000" else
			"1111110010010110" when input = "0000000011010001" else
			"1111110010011110" when input = "0000000011010010" else
			"1111110010100111" when input = "0000000011010011" else
			"1111110010110000" when input = "0000000011010100" else
			"1111110010111010" when input = "0000000011010101" else
			"1111110011000011" when input = "0000000011010110" else
			"1111110011001101" when input = "0000000011010111" else
			"1111110011010111" when input = "0000000011011000" else
			"1111110011100010" when input = "0000000011011001" else
			"1111110011101100" when input = "0000000011011010" else
			"1111110011110111" when input = "0000000011011011" else
			"1111110100000010" when input = "0000000011011100" else
			"1111110100001110" when input = "0000000011011101" else
			"1111110100011001" when input = "0000000011011110" else
			"1111110100100101" when input = "0000000011011111" else
			"1111110100110001" when input = "0000000011100000" else
			"1111110100111101" when input = "0000000011100001" else
			"1111110101001010" when input = "0000000011100010" else
			"1111110101010110" when input = "0000000011100011" else
			"1111110101100011" when input = "0000000011100100" else
			"1111110101110000" when input = "0000000011100101" else
			"1111110101111110" when input = "0000000011100110" else
			"1111110110001011" when input = "0000000011100111" else
			"1111110110011001" when input = "0000000011101000" else
			"1111110110100111" when input = "0000000011101001" else
			"1111110110110101" when input = "0000000011101010" else
			"1111110111000011" when input = "0000000011101011" else
			"1111110111010001" when input = "0000000011101100" else
			"1111110111100000" when input = "0000000011101101" else
			"1111110111101110" when input = "0000000011101110" else
			"1111110111111101" when input = "0000000011101111" else
			"1111111000001100" when input = "0000000011110000" else
			"1111111000011100" when input = "0000000011110001" else
			"1111111000101011" when input = "0000000011110010" else
			"1111111000111010" when input = "0000000011110011" else
			"1111111001001010" when input = "0000000011110100" else
			"1111111001011010" when input = "0000000011110101" else
			"1111111001101010" when input = "0000000011110110" else
			"1111111001111010" when input = "0000000011110111" else
			"1111111010001010" when input = "0000000011111000" else
			"1111111010011010" when input = "0000000011111001" else
			"1111111010101010" when input = "0000000011111010" else
			"1111111010111011" when input = "0000000011111011" else
			"1111111011001011" when input = "0000000011111100" else
			"1111111011011100" when input = "0000000011111101" else
			"1111111011101101" when input = "0000000011111110" else
			"1111111011111110" when input = "0000000011111111" else
			"1111111100001110" when input = "0000000100000000" else
			"1111111100011111" when input = "0000000100000001" else
			"1111111100110000" when input = "0000000100000010" else
			"1111111101000010" when input = "0000000100000011" else
			"1111111101010011" when input = "0000000100000100" else
			"1111111101100100" when input = "0000000100000101" else
			"1111111101110101" when input = "0000000100000110" else
			"1111111110000110" when input = "0000000100000111" else
			"1111111110011000" when input = "0000000100001000" else
			"1111111110101001" when input = "0000000100001001" else
			"1111111110111011" when input = "0000000100001010" else
			"1111111111001100" when input = "0000000100001011" else
			"1111111111011101" when input = "0000000100001100" else
			"1111111111101111" when input = "0000000100001101" else
			"0000000000000000" when input = "0000000100001110" else
			"0000000000010001" when input = "0000000100001111" else
			"0000000000100010" when input = "0000000100010000" else
			"0000000000110100" when input = "0000000100010001" else
			"0000000001000101" when input = "0000000100010010" else
			"0000000001010111" when input = "0000000100010011" else
			"0000000001101000" when input = "0000000100010100" else
			"0000000001111001" when input = "0000000100010101" else
			"0000000010001011" when input = "0000000100010110" else
			"0000000010011100" when input = "0000000100010111" else
			"0000000010101101" when input = "0000000100011000" else
			"0000000010111110" when input = "0000000100011001" else
			"0000000011001111" when input = "0000000100011010" else
			"0000000011100000" when input = "0000000100011011" else
			"0000000011110001" when input = "0000000100011100" else
			"0000000100000010" when input = "0000000100011101" else
			"0000000100010011" when input = "0000000100011110" else
			"0000000100100100" when input = "0000000100011111" else
			"0000000100110100" when input = "0000000100100000" else
			"0000000101000101" when input = "0000000100100001" else
			"0000000101010101" when input = "0000000100100010" else
			"0000000101100110" when input = "0000000100100011" else
			"0000000101110110" when input = "0000000100100100" else
			"0000000110000110" when input = "0000000100100101" else
			"0000000110010110" when input = "0000000100100110" else
			"0000000110100110" when input = "0000000100100111" else
			"0000000110110110" when input = "0000000100101000" else
			"0000000111000101" when input = "0000000100101001" else
			"0000000111010101" when input = "0000000100101010" else
			"0000000111100100" when input = "0000000100101011" else
			"0000000111110011" when input = "0000000100101100" else
			"0000001000000010" when input = "0000000100101101" else
			"0000001000010001" when input = "0000000100101110" else
			"0000001000100000" when input = "0000000100101111" else
			"0000001000101111" when input = "0000000100110000" else
			"0000001000111101" when input = "0000000100110001" else
			"0000001001001011" when input = "0000000100110010" else
			"0000001001011001" when input = "0000000100110011" else
			"0000001001100111" when input = "0000000100110100" else
			"0000001001110101" when input = "0000000100110101" else
			"0000001010000010" when input = "0000000100110110" else
			"0000001010001111" when input = "0000000100110111" else
			"0000001010011101" when input = "0000000100111000" else
			"0000001010101001" when input = "0000000100111001" else
			"0000001010110110" when input = "0000000100111010" else
			"0000001011000010" when input = "0000000100111011" else
			"0000001011001111" when input = "0000000100111100" else
			"0000001011011011" when input = "0000000100111101" else
			"0000001011100111" when input = "0000000100111110" else
			"0000001011110010" when input = "0000000100111111" else
			"0000001011111101" when input = "0000000101000000" else
			"0000001100001001" when input = "0000000101000001" else
			"0000001100010011" when input = "0000000101000010" else
			"0000001100011110" when input = "0000000101000011" else
			"0000001100101000" when input = "0000000101000100" else
			"0000001100110011" when input = "0000000101000101" else
			"0000001100111100" when input = "0000000101000110" else
			"0000001101000110" when input = "0000000101000111" else
			"0000001101001111" when input = "0000000101001000" else
			"0000001101011001" when input = "0000000101001001" else
			"0000001101100001" when input = "0000000101001010" else
			"0000001101101010" when input = "0000000101001011" else
			"0000001101110010" when input = "0000000101001100" else
			"0000001101111010" when input = "0000000101001101" else
			"0000001110000010" when input = "0000000101001110" else
			"0000001110001010" when input = "0000000101001111" else
			"0000001110010001" when input = "0000000101010000" else
			"0000001110011000" when input = "0000000101010001" else
			"0000001110011111" when input = "0000000101010010" else
			"0000001110100101" when input = "0000000101010011" else
			"0000001110101011" when input = "0000000101010100" else
			"0000001110110001" when input = "0000000101010101" else
			"0000001110110111" when input = "0000000101010110" else
			"0000001110111100" when input = "0000000101010111" else
			"0000001111000001" when input = "0000000101011000" else
			"0000001111000101" when input = "0000000101011001" else
			"0000001111001010" when input = "0000000101011010" else
			"0000001111001110" when input = "0000000101011011" else
			"0000001111010010" when input = "0000000101011100" else
			"0000001111010101" when input = "0000000101011101" else
			"0000001111011000" when input = "0000000101011110" else
			"0000001111011011" when input = "0000000101011111" else
			"0000001111011110" when input = "0000000101100000" else
			"0000001111100000" when input = "0000000101100001" else
			"0000001111100010" when input = "0000000101100010" else
			"0000001111100100" when input = "0000000101100011" else
			"0000001111100101" when input = "0000000101100100" else
			"0000001111100110" when input = "0000000101100101" else
			"0000001111100111" when input = "0000000101100110" else
			"0000001111100111" when input = "0000000101100111" else
			"0000001111100111" when input = "0000000101101000" else
			"XXXXXXXXXXXXXXXX";
end architecture ;
