library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity sqrt_co is
	port (
	input : in std_logic_vector(15 DOWNTO 0);
	output : out std_logic_vector(15 DOWNTO 0)
	);
end sqrt_co;

architecture rtl of sqrt_co is
begin
	output <=
			"0000000000000000" when input <= "0000000000000001" else
			"0000000000000010" when input <= "0000000000000100" else
			"0000000000000011" when input <= "0000000000001001" else
			"0000000000000100" when input <= "0000000000010000" else
			"0000000000000101" when input <= "0000000000011001" else
			"0000000000000110" when input <= "0000000000100100" else
			"0000000000000111" when input <= "0000000000110001" else
			"0000000000001000" when input <= "0000000001000000" else
			"0000000000001001" when input <= "0000000001010001" else
			"0000000000001010" when input <= "0000000001100100" else
			"0000000000001011" when input <= "0000000001111001" else
			"0000000000001100" when input <= "0000000010010000" else
			"0000000000001101" when input <= "0000000010101001" else
			"0000000000001110" when input <= "0000000011000100" else
			"0000000000001111" when input <= "0000000011100001" else
			"0000000000010000" when input <= "0000000100000000" else
			"0000000000010001" when input <= "0000000100100001" else
			"0000000000010010" when input <= "0000000101000100" else
			"0000000000010011" when input <= "0000000101101001" else
			"0000000000010100" when input <= "0000000110010000" else
			"0000000000010101" when input <= "0000000110111001" else
			"0000000000010110" when input <= "0000000111100100" else
			"0000000000010111" when input <= "0000001000010001" else
			"0000000000011000" when input <= "0000001001000000" else
			"0000000000011001" when input <= "0000001001110001" else
			"0000000000011010" when input <= "0000001010100100" else
			"0000000000011011" when input <= "0000001011011001" else
			"0000000000011100" when input <= "0000001100010000" else
			"0000000000011101" when input <= "0000001101001001" else
			"0000000000011110" when input <= "0000001110000100" else
			"0000000000011111" when input <= "0000001111000001" else
			"0000000000100000" when input <= "0000010000000000" else
			"0000000000100001" when input <= "0000010001000001" else
			"0000000000100010" when input <= "0000010010000100" else
			"0000000000100011" when input <= "0000010011001001" else
			"0000000000100100" when input <= "0000010100010000" else
			"0000000000100101" when input <= "0000010101011001" else
			"0000000000100110" when input <= "0000010110100100" else
			"0000000000100111" when input <= "0000010111110001" else
			"0000000000101000" when input <= "0000011001000000" else
			"0000000000101001" when input <= "0000011010010001" else
			"0000000000101010" when input <= "0000011011100100" else
			"0000000000101011" when input <= "0000011100111001" else
			"0000000000101100" when input <= "0000011110010000" else
			"0000000000101101" when input <= "0000011111101001" else
			"0000000000101110" when input <= "0000100001000100" else
			"0000000000101111" when input <= "0000100010100001" else
			"0000000000110000" when input <= "0000100100000000" else
			"0000000000110001" when input <= "0000100101100001" else
			"0000000000110010" when input <= "0000100111000100" else
			"0000000000110011" when input <= "0000101000101001" else
			"0000000000110100" when input <= "0000101010010000" else
			"0000000000110101" when input <= "0000101011111001" else
			"0000000000110110" when input <= "0000101101100100" else
			"0000000000110111" when input <= "0000101111010001" else
			"0000000000111000" when input <= "0000110001000000" else
			"0000000000111001" when input <= "0000110010110001" else
			"0000000000111010" when input <= "0000110100100100" else
			"0000000000111011" when input <= "0000110110011001" else
			"0000000000111100" when input <= "0000111000010000" else
			"0000000000111101" when input <= "0000111010001001" else
			"0000000000111110" when input <= "0000111100000100" else
			"0000000000111111" when input <= "0000111110000001" else
			"0000000001000000" when input <= "0001000000000000" else
			"0000000001000001" when input <= "0001000010000001" else
			"0000000001000010" when input <= "0001000100000100" else
			"0000000001000011" when input <= "0001000110001001" else
			"0000000001000100" when input <= "0001001000010000" else
			"0000000001000101" when input <= "0001001010011001" else
			"0000000001000110" when input <= "0001001100100100" else
			"0000000001000111" when input <= "0001001110110001" else
			"0000000001001000" when input <= "0001010001000000" else
			"0000000001001001" when input <= "0001010011010001" else
			"0000000001001010" when input <= "0001010101100100" else
			"0000000001001011" when input <= "0001010111111001" else
			"0000000001001100" when input <= "0001011010010000" else
			"0000000001001101" when input <= "0001011100101001" else
			"0000000001001110" when input <= "0001011111000100" else
			"0000000001001111" when input <= "0001100001100001" else
			"0000000001010000" when input <= "0001100100000000" else
			"0000000001010001" when input <= "0001100110100001" else
			"0000000001010010" when input <= "0001101001000100" else
			"0000000001010011" when input <= "0001101011101001" else
			"0000000001010100" when input <= "0001101110010000" else
			"0000000001010101" when input <= "0001110000111001" else
			"0000000001010110" when input <= "0001110011100100" else
			"0000000001010111" when input <= "0001110110010001" else
			"0000000001011000" when input <= "0001111001000000" else
			"0000000001011001" when input <= "0001111011110001" else
			"0000000001011010" when input <= "0001111110100100" else
			"0000000001011011" when input <= "0010000001011001" else
			"0000000001011100" when input <= "0010000100010000" else
			"0000000001011101" when input <= "0010000111001001" else
			"0000000001011110" when input <= "0010001010000100" else
			"0000000001011111" when input <= "0010001101000001" else
			"0000000001100000" when input <= "0010010000000000" else
			"0000000001100001" when input <= "0010010011000001" else
			"0000000001100010" when input <= "0010010110000100" else
			"0000000001100011" when input <= "0010011001001001" else
			"0000000001100100" when input <= "0010011100010000" else
			"0000000001100101" when input <= "0010011111011001" else
			"0000000001100110" when input <= "0010100010100100" else
			"0000000001100111" when input <= "0010100101110001" else
			"0000000001101000" when input <= "0010101001000000" else
			"0000000001101001" when input <= "0010101100010001" else
			"0000000001101010" when input <= "0010101111100100" else
			"0000000001101011" when input <= "0010110010111001" else
			"0000000001101100" when input <= "0010110110010000" else
			"0000000001101101" when input <= "0010111001101001" else
			"0000000001101110" when input <= "0010111101000100" else
			"0000000001101111" when input <= "0011000000100001" else
			"0000000001110000" when input <= "0011000100000000" else
			"0000000001110001" when input <= "0011000111100001" else
			"0000000001110010" when input <= "0011001011000100" else
			"0000000001110011" when input <= "0011001110101001" else
			"0000000001110100" when input <= "0011010010010000" else
			"0000000001110101" when input <= "0011010101111001" else
			"0000000001110110" when input <= "0011011001100100" else
			"0000000001110111" when input <= "0011011101010001" else
			"0000000001111000" when input <= "0011100001000000" else
			"0000000001111001" when input <= "0011100100110001" else
			"0000000001111010" when input <= "0011101000100100" else
			"0000000001111011" when input <= "0011101100011001" else
			"0000000001111100" when input <= "0011110000010000" else
			"0000000001111101" when input <= "0011110100001001" else
			"0000000001111110" when input <= "0011111000000100" else
			"0000000001111111" when input <= "0011111100000001" else
			"0000000010000000" when input <= "0100000000000000" else
			"0000000010000001" when input <= "0100000100000001" else
			"0000000010000010" when input <= "0100001000000100" else
			"0000000010000011" when input <= "0100001100001001" else
			"0000000010000100" when input <= "0100010000010000" else
			"0000000010000101" when input <= "0100010100011001" else
			"0000000010000110" when input <= "0100011000100100" else
			"0000000010000111" when input <= "0100011100110001" else
			"0000000010001000" when input <= "0100100001000000" else
			"0000000010001001" when input <= "0100100101010001" else
			"0000000010001010" when input <= "0100101001100100" else
			"0000000010001011" when input <= "0100101101111001" else
			"0000000010001100" when input <= "0100110010010000" else
			"0000000010001101" when input <= "0100110110101001" else
			"0000000010001110" when input <= "0100111011000100" else
			"0000000010001111" when input <= "0100111111100001" else
			"0000000010010000" when input <= "0101000100000000" else
			"0000000010010001" when input <= "0101001000100001" else
			"0000000010010010" when input <= "0101001101000100" else
			"0000000010010011" when input <= "0101010001101001" else
			"0000000010010100" when input <= "0101010110010000" else
			"0000000010010101" when input <= "0101011010111001" else
			"0000000010010110" when input <= "0101011111100100" else
			"0000000010010111" when input <= "0101100100010001" else
			"0000000010011000" when input <= "0101101001000000" else
			"0000000010011001" when input <= "0101101101110001" else
			"0000000010011010" when input <= "0101110010100100" else
			"0000000010011011" when input <= "0101110111011001" else
			"0000000010011100" when input <= "0101111100010000" else
			"0000000010011101" when input <= "0110000001001001" else
			"0000000010011110" when input <= "0110000110000100" else
			"0000000010011111" when input <= "0110001011000001" else
			"0000000010100000" when input <= "0110010000000000" else
			"0000000010100001" when input <= "0110010101000001" else
			"0000000010100010" when input <= "0110011010000100" else
			"0000000010100011" when input <= "0110011111001001" else
			"0000000010100100" when input <= "0110100100010000" else
			"0000000010100101" when input <= "0110101001011001" else
			"0000000010100110" when input <= "0110101110100100" else
			"0000000010100111" when input <= "0110110011110001" else
			"0000000010101000" when input <= "0110111001000000" else
			"0000000010101001" when input <= "0110111110010001" else
			"0000000010101010" when input <= "0111000011100100" else
			"0000000010101011" when input <= "0111001000111001" else
			"0000000010101100" when input <= "0111001110010000" else
			"0000000010101101" when input <= "0111010011101001" else
			"0000000010101110" when input <= "0111011001000100" else
			"0000000010101111" when input <= "0111011110100001" else
			"0000000010110000" when input <= "0111100100000000" else
			"0000000010110001" when input <= "0111101001100001" else
			"0000000010110010" when input <= "0111101111000100" else
			"0000000010110011" when input <= "0111110100101001" else
			"0000000010110100" when input <= "0111111010010000" else
			"0000000010110101" when input <= "0111111111111001" else
			"XXXXXXXXXXXXXXXX";
end architecture ;
